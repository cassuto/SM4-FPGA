
module sbox_8b(
   input CLK_i,
   input [7:0] X_i,
   output reg [7:0] Y_o
);

   /* sbox ROM */
   always @(posedge CLK_i) begin
      case (X_i)
         8'h00: Y_o <= 8'hD6;
         8'h01: Y_o <= 8'h90;
         8'h02: Y_o <= 8'hE9;
         8'h03: Y_o <= 8'hFE;
         8'h04: Y_o <= 8'hCC;
         8'h05: Y_o <= 8'hE1;
         8'h06: Y_o <= 8'h3D;
         8'h07: Y_o <= 8'hB7;
         8'h08: Y_o <= 8'h16;
         8'h09: Y_o <= 8'hB6;
         8'h0A: Y_o <= 8'h14;
         8'h0B: Y_o <= 8'hC2;
         8'h0C: Y_o <= 8'h28;
         8'h0D: Y_o <= 8'hFB;
         8'h0E: Y_o <= 8'h2C;
         8'h0F: Y_o <= 8'h05;
         8'h10: Y_o <= 8'h2B;
         8'h11: Y_o <= 8'h67;
         8'h12: Y_o <= 8'h9A;
         8'h13: Y_o <= 8'h76;
         8'h14: Y_o <= 8'h2A;
         8'h15: Y_o <= 8'hBE;
         8'h16: Y_o <= 8'h04;
         8'h17: Y_o <= 8'hC3;
         8'h18: Y_o <= 8'hAA;
         8'h19: Y_o <= 8'h44;
         8'h1A: Y_o <= 8'h13;
         8'h1B: Y_o <= 8'h26;
         8'h1C: Y_o <= 8'h49;
         8'h1D: Y_o <= 8'h86;
         8'h1E: Y_o <= 8'h06;
         8'h1F: Y_o <= 8'h99;
         8'h20: Y_o <= 8'h9C;
         8'h21: Y_o <= 8'h42;
         8'h22: Y_o <= 8'h50;
         8'h23: Y_o <= 8'hF4;
         8'h24: Y_o <= 8'h91;
         8'h25: Y_o <= 8'hEF;
         8'h26: Y_o <= 8'h98;
         8'h27: Y_o <= 8'h7A;
         8'h28: Y_o <= 8'h33;
         8'h29: Y_o <= 8'h54;
         8'h2A: Y_o <= 8'h0B;
         8'h2B: Y_o <= 8'h43;
         8'h2C: Y_o <= 8'hED;
         8'h2D: Y_o <= 8'hCF;
         8'h2E: Y_o <= 8'hAC;
         8'h2F: Y_o <= 8'h62;
         8'h30: Y_o <= 8'hE4;
         8'h31: Y_o <= 8'hB3;
         8'h32: Y_o <= 8'h1C;
         8'h33: Y_o <= 8'hA9;
         8'h34: Y_o <= 8'hC9;
         8'h35: Y_o <= 8'h08;
         8'h36: Y_o <= 8'hE8;
         8'h37: Y_o <= 8'h95;
         8'h38: Y_o <= 8'h80;
         8'h39: Y_o <= 8'hDF;
         8'h3A: Y_o <= 8'h94;
         8'h3B: Y_o <= 8'hFA;
         8'h3C: Y_o <= 8'h75;
         8'h3D: Y_o <= 8'h8F;
         8'h3E: Y_o <= 8'h3F;
         8'h3F: Y_o <= 8'hA6;
         8'h40: Y_o <= 8'h47;
         8'h41: Y_o <= 8'h07;
         8'h42: Y_o <= 8'hA7;
         8'h43: Y_o <= 8'hFC;
         8'h44: Y_o <= 8'hF3;
         8'h45: Y_o <= 8'h73;
         8'h46: Y_o <= 8'h17;
         8'h47: Y_o <= 8'hBA;
         8'h48: Y_o <= 8'h83;
         8'h49: Y_o <= 8'h59;
         8'h4A: Y_o <= 8'h3C;
         8'h4B: Y_o <= 8'h19;
         8'h4C: Y_o <= 8'hE6;
         8'h4D: Y_o <= 8'h85;
         8'h4E: Y_o <= 8'h4F;
         8'h4F: Y_o <= 8'hA8;
         8'h50: Y_o <= 8'h68;
         8'h51: Y_o <= 8'h6B;
         8'h52: Y_o <= 8'h81;
         8'h53: Y_o <= 8'hB2;
         8'h54: Y_o <= 8'h71;
         8'h55: Y_o <= 8'h64;
         8'h56: Y_o <= 8'hDA;
         8'h57: Y_o <= 8'h8B;
         8'h58: Y_o <= 8'hF8;
         8'h59: Y_o <= 8'hEB;
         8'h5A: Y_o <= 8'h0F;
         8'h5B: Y_o <= 8'h4B;
         8'h5C: Y_o <= 8'h70;
         8'h5D: Y_o <= 8'h56;
         8'h5E: Y_o <= 8'h9D;
         8'h5F: Y_o <= 8'h35;
         8'h60: Y_o <= 8'h1E;
         8'h61: Y_o <= 8'h24;
         8'h62: Y_o <= 8'h0E;
         8'h63: Y_o <= 8'h5E;
         8'h64: Y_o <= 8'h63;
         8'h65: Y_o <= 8'h58;
         8'h66: Y_o <= 8'hD1;
         8'h67: Y_o <= 8'hA2;
         8'h68: Y_o <= 8'h25;
         8'h69: Y_o <= 8'h22;
         8'h6A: Y_o <= 8'h7C;
         8'h6B: Y_o <= 8'h3B;
         8'h6C: Y_o <= 8'h01;
         8'h6D: Y_o <= 8'h21;
         8'h6E: Y_o <= 8'h78;
         8'h6F: Y_o <= 8'h87;
         8'h70: Y_o <= 8'hD4;
         8'h71: Y_o <= 8'h00;
         8'h72: Y_o <= 8'h46;
         8'h73: Y_o <= 8'h57;
         8'h74: Y_o <= 8'h9F;
         8'h75: Y_o <= 8'hD3;
         8'h76: Y_o <= 8'h27;
         8'h77: Y_o <= 8'h52;
         8'h78: Y_o <= 8'h4C;
         8'h79: Y_o <= 8'h36;
         8'h7A: Y_o <= 8'h02;
         8'h7B: Y_o <= 8'hE7;
         8'h7C: Y_o <= 8'hA0;
         8'h7D: Y_o <= 8'hC4;
         8'h7E: Y_o <= 8'hC8;
         8'h7F: Y_o <= 8'h9E;
         8'h80: Y_o <= 8'hEA;
         8'h81: Y_o <= 8'hBF;
         8'h82: Y_o <= 8'h8A;
         8'h83: Y_o <= 8'hD2;
         8'h84: Y_o <= 8'h40;
         8'h85: Y_o <= 8'hC7;
         8'h86: Y_o <= 8'h38;
         8'h87: Y_o <= 8'hB5;
         8'h88: Y_o <= 8'hA3;
         8'h89: Y_o <= 8'hF7;
         8'h8A: Y_o <= 8'hF2;
         8'h8B: Y_o <= 8'hCE;
         8'h8C: Y_o <= 8'hF9;
         8'h8D: Y_o <= 8'h61;
         8'h8E: Y_o <= 8'h15;
         8'h8F: Y_o <= 8'hA1;
         8'h90: Y_o <= 8'hE0;
         8'h91: Y_o <= 8'hAE;
         8'h92: Y_o <= 8'h5D;
         8'h93: Y_o <= 8'hA4;
         8'h94: Y_o <= 8'h9B;
         8'h95: Y_o <= 8'h34;
         8'h96: Y_o <= 8'h1A;
         8'h97: Y_o <= 8'h55;
         8'h98: Y_o <= 8'hAD;
         8'h99: Y_o <= 8'h93;
         8'h9A: Y_o <= 8'h32;
         8'h9B: Y_o <= 8'h30;
         8'h9C: Y_o <= 8'hF5;
         8'h9D: Y_o <= 8'h8C;
         8'h9E: Y_o <= 8'hB1;
         8'h9F: Y_o <= 8'hE3;
         8'hA0: Y_o <= 8'h1D;
         8'hA1: Y_o <= 8'hF6;
         8'hA2: Y_o <= 8'hE2;
         8'hA3: Y_o <= 8'h2E;
         8'hA4: Y_o <= 8'h82;
         8'hA5: Y_o <= 8'h66;
         8'hA6: Y_o <= 8'hCA;
         8'hA7: Y_o <= 8'h60;
         8'hA8: Y_o <= 8'hC0;
         8'hA9: Y_o <= 8'h29;
         8'hAA: Y_o <= 8'h23;
         8'hAB: Y_o <= 8'hAB;
         8'hAC: Y_o <= 8'h0D;
         8'hAD: Y_o <= 8'h53;
         8'hAE: Y_o <= 8'h4E;
         8'hAF: Y_o <= 8'h6F;
         8'hB0: Y_o <= 8'hD5;
         8'hB1: Y_o <= 8'hDB;
         8'hB2: Y_o <= 8'h37;
         8'hB3: Y_o <= 8'h45;
         8'hB4: Y_o <= 8'hDE;
         8'hB5: Y_o <= 8'hFD;
         8'hB6: Y_o <= 8'h8E;
         8'hB7: Y_o <= 8'h2F;
         8'hB8: Y_o <= 8'h03;
         8'hB9: Y_o <= 8'hFF;
         8'hBA: Y_o <= 8'h6A;
         8'hBB: Y_o <= 8'h72;
         8'hBC: Y_o <= 8'h6D;
         8'hBD: Y_o <= 8'h6C;
         8'hBE: Y_o <= 8'h5B;
         8'hBF: Y_o <= 8'h51;
         8'hC0: Y_o <= 8'h8D;
         8'hC1: Y_o <= 8'h1B;
         8'hC2: Y_o <= 8'hAF;
         8'hC3: Y_o <= 8'h92;
         8'hC4: Y_o <= 8'hBB;
         8'hC5: Y_o <= 8'hDD;
         8'hC6: Y_o <= 8'hBC;
         8'hC7: Y_o <= 8'h7F;
         8'hC8: Y_o <= 8'h11;
         8'hC9: Y_o <= 8'hD9;
         8'hCA: Y_o <= 8'h5C;
         8'hCB: Y_o <= 8'h41;
         8'hCC: Y_o <= 8'h1F;
         8'hCD: Y_o <= 8'h10;
         8'hCE: Y_o <= 8'h5A;
         8'hCF: Y_o <= 8'hD8;
         8'hD0: Y_o <= 8'h0A;
         8'hD1: Y_o <= 8'hC1;
         8'hD2: Y_o <= 8'h31;
         8'hD3: Y_o <= 8'h88;
         8'hD4: Y_o <= 8'hA5;
         8'hD5: Y_o <= 8'hCD;
         8'hD6: Y_o <= 8'h7B;
         8'hD7: Y_o <= 8'hBD;
         8'hD8: Y_o <= 8'h2D;
         8'hD9: Y_o <= 8'h74;
         8'hDA: Y_o <= 8'hD0;
         8'hDB: Y_o <= 8'h12;
         8'hDC: Y_o <= 8'hB8;
         8'hDD: Y_o <= 8'hE5;
         8'hDE: Y_o <= 8'hB4;
         8'hDF: Y_o <= 8'hB0;
         8'hE0: Y_o <= 8'h89;
         8'hE1: Y_o <= 8'h69;
         8'hE2: Y_o <= 8'h97;
         8'hE3: Y_o <= 8'h4A;
         8'hE4: Y_o <= 8'h0C;
         8'hE5: Y_o <= 8'h96;
         8'hE6: Y_o <= 8'h77;
         8'hE7: Y_o <= 8'h7E;
         8'hE8: Y_o <= 8'h65;
         8'hE9: Y_o <= 8'hB9;
         8'hEA: Y_o <= 8'hF1;
         8'hEB: Y_o <= 8'h09;
         8'hEC: Y_o <= 8'hC5;
         8'hED: Y_o <= 8'h6E;
         8'hEE: Y_o <= 8'hC6;
         8'hEF: Y_o <= 8'h84;
         8'hF0: Y_o <= 8'h18;
         8'hF1: Y_o <= 8'hF0;
         8'hF2: Y_o <= 8'h7D;
         8'hF3: Y_o <= 8'hEC;
         8'hF4: Y_o <= 8'h3A;
         8'hF5: Y_o <= 8'hDC;
         8'hF6: Y_o <= 8'h4D;
         8'hF7: Y_o <= 8'h20;
         8'hF8: Y_o <= 8'h79;
         8'hF9: Y_o <= 8'hEE;
         8'hFA: Y_o <= 8'h5F;
         8'hFB: Y_o <= 8'h3E;
         8'hFC: Y_o <= 8'hD7;
         8'hFD: Y_o <= 8'hCB;
         8'hFE: Y_o <= 8'h39;
         8'hFF: Y_o <= 8'h48;
      endcase
   end

endmodule
